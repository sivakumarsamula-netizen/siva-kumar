class tb;
	int a,b;

	initial begin
		
		$display("siva kumar samula");
		$display("hiiiiiii");

	end

endclass
